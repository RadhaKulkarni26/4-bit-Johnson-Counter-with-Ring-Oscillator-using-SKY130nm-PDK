* /home/radhadk260501/eSim-Workspace/Radha_Johnson_Counter/Radha_Johnson_Counter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 08 Oct 2022 03:26:00 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ counter_module		
U3  clk T Net-_U2-Pad1_ Net-_U2-Pad2_ adc_bridge_2		
U4  Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ A B C D dac_bridge_4		
SC7  Net-_SC1-Pad2_ clk Net-_SC1-Pad3_ sky130_fd_pr__res_generic_nd		
SC8  clk GND Net-_SC1-Pad3_ sky130_fd_pr__res_generic_nd		
v2  Net-_SC1-Pad3_ GND DC		
scmode1  SKY130mode		
U5  clk plot_v1		
U6  A plot_v1		
U7  B plot_v1		
U8  C plot_v1		
U9  D plot_v1		
SC2  Net-_SC1-Pad1_ Net-_SC1-Pad2_ GND GND sky130_fd_pr__nfet_01v8_lvt		
SC4  Net-_SC3-Pad1_ Net-_SC1-Pad1_ GND GND sky130_fd_pr__nfet_01v8_lvt		
SC6  Net-_SC1-Pad2_ Net-_SC3-Pad1_ GND GND sky130_fd_pr__nfet_01v8_lvt		
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8_lvt		
SC3  Net-_SC3-Pad1_ Net-_SC1-Pad1_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8_lvt		
SC5  Net-_SC1-Pad2_ Net-_SC3-Pad1_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8_lvt		
U1  T plot_v1		
v1  T GND pulse		

.end
